--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:05:11 05/04/2019
-- Design Name:   
-- Module Name:   /home/ajd12342/CS-226-Project/classify_tb.vhd
-- Project Name:  classify
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: classify_packet
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY classify_tb IS
END classify_tb;
 
ARCHITECTURE behavior OF classify_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT classify_packet
    PORT(
         iData_av : IN  std_logic_vector(31 downto 0);
         iRd_Data : OUT  std_logic_vector(31 downto 0);
         iData0 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData1 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData2 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData3 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData4 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData5 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData6 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData7 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData8 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData9 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData10 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData11 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData12 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData13 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData14 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData15 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData16 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData17 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData18 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData19 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData20 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData21 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData22 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData23 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData24 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData25 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData26 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData27 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData28 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData29 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData30 : in  STD_LOGIC_VECTOR (143 downto 0);
    		  iData31 : in  STD_LOGIC_VECTOR (143 downto 0);
         oData_av : OUT  std_logic;
         oData_rd : IN  std_logic;
         oData : OUT  std_logic_vector(143 downto 0);
         MAC : IN  std_logic_vector(47 downto 0);
         valid_in : IN  std_logic;
         valid_out : OUT  std_logic;
         Opcode : OUT  std_logic_vector(2 downto 0);
         Rd_opcode : IN  std_logic;
         Input_port : OUT  std_logic_vector(4 downto 0);
         Port_mask : OUT  std_logic_vector(31 downto 0);
         Edge_ports : INOUT  std_logic_vector(31 downto 0);
         Core_Ports : INOUT  std_logic_vector(31 downto 0);
         gport : OUT  std_logic_vector(31 downto 0);
         ostatus : OUT  std_logic_vector(1 downto 0);
         oreadstatus : OUT  std_logic_vector(3 downto 0);
         debug : INOUT  std_logic_vector(15 downto 0);
         hoppointer_o : OUT  std_logic_vector(15 downto 0);
         pkt0_0 : OUT  std_logic_vector(144 downto 0);
         pkt1_0 : OUT  std_logic_vector(144 downto 0);
         pkt2_0 : OUT  std_logic_vector(144 downto 0);
         pkt3_0 : OUT  std_logic_vector(144 downto 0);
         pkt4_0 : OUT  std_logic_vector(144 downto 0);
         counter_o : OUT  std_logic_vector(23 downto 0);
         ethertype_o : OUT  std_logic_vector(15 downto 0);
         ethervalue_o : OUT  std_logic_vector(15 downto 0);
         counter_index : OUT  integer range 0 to 15;
         grantportint_o : OUT  integer range 1 to 32;
         addlpointer_o : OUT  integer range 0 to 479;
         addrpointer_o : OUT  integer range 0 to 479;
         ready2push_o : OUT  std_logic;
         dropped_o : OUT  std_logic;
         isfull_o : OUT  std_logic;
         clk : IN  std_logic;
         rst : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal iData_av : std_logic_vector(31 downto 0) := (others => '0');
	signal iData0 :  STD_LOGIC_VECTOR (143 downto 0);
  signal iData1 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData2 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData3 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData4 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData5 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData6 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData7 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData8 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData9 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData10 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData11 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData12 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData13 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData14 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData15 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData16 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData17 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData18 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData19 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData20 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData21 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData22 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData23 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData24 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData25 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData26 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData27 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData28 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData29 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData30 : STD_LOGIC_VECTOR (143 downto 0);
  signal iData31 : STD_LOGIC_VECTOR (143 downto 0);
   signal oData_rd : std_logic := '0';
   signal MAC : std_logic_vector(47 downto 0) := (others => '0');
   signal valid_in : std_logic := '0';
   signal Rd_opcode : std_logic := '0';
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';

	--BiDirs
   signal Edge_ports : std_logic_vector(31 downto 0);
   signal Core_Ports : std_logic_vector(31 downto 0);
   signal debug : std_logic_vector(15 downto 0);

 	--Outputs
   signal iRd_Data : std_logic_vector(31 downto 0);
   signal oData_av : std_logic;
   signal oData : std_logic_vector(143 downto 0);
   signal valid_out : std_logic;
   signal Opcode : std_logic_vector(2 downto 0);
   signal Input_port : std_logic_vector(4 downto 0);
   signal Port_mask : std_logic_vector(31 downto 0);
   signal gport : std_logic_vector(31 downto 0);
   signal ostatus : std_logic_vector(1 downto 0);
   signal oreadstatus : std_logic_vector(3 downto 0);
   signal hoppointer_o : std_logic_vector(15 downto 0);
   signal pkt0_0 : std_logic_vector(144 downto 0);
   signal pkt1_0 : std_logic_vector(144 downto 0);
   signal pkt2_0 : std_logic_vector(144 downto 0);
   signal pkt3_0 : std_logic_vector(144 downto 0);
   signal pkt4_0 : std_logic_vector(144 downto 0);
   signal counter_o : std_logic_vector(23 downto 0);
   signal ethertype_o : std_logic_vector(15 downto 0);
   signal ethervalue_o : std_logic_vector(15 downto 0);
   signal counter_index : integer range 0 to 15;
   signal grantportint_o : integer range 1 to 32;
   signal addlpointer_o : integer range 0 to 479;
   signal addrpointer_o : integer range 0 to 479;
   signal ready2push_o : std_logic;
   signal dropped_o : std_logic;
   signal isfull_o : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: classify_packet PORT MAP (
          iData_av => iData_av,
          iRd_Data => iRd_Data,
          iData0 => iData0,
iData1 => iData1,
iData2 => iData2,
iData3 => iData3,
iData4 => iData4,
iData5 => iData5,
iData6 => iData6,
iData7 => iData7,
iData8 => iData8,
iData9 => iData9,
iData10 => iData10,
iData11 => iData11,
iData12 => iData12,
iData13 => iData13,
iData14 => iData14,
iData15 => iData15,
iData16 => iData16,
iData17 => iData17,
iData18 => iData18,
iData19 => iData19,
iData20 => iData20,
iData21 => iData21,
iData22 => iData22,
iData23 => iData23,
iData24 => iData24,
iData25 => iData25,
iData26 => iData26,
iData27 => iData27,
iData28 => iData28,
iData29 => iData29,
iData30 => iData30,
iData31 => iData31,

          oData_av => oData_av,
          oData_rd => oData_rd,
          oData => oData,
          MAC => MAC,
          valid_in => valid_in,
          valid_out => valid_out,
          Opcode => Opcode,
          Rd_opcode => Rd_opcode,
          Input_port => Input_port,
          Port_mask => Port_mask,
          Edge_ports => Edge_ports,
          Core_Ports => Core_Ports,
          gport => gport,
          ostatus => ostatus,
          oreadstatus => oreadstatus,
          debug => debug,
          hoppointer_o => hoppointer_o,
          pkt0_0 => pkt0_0,
          pkt1_0 => pkt1_0,
          pkt2_0 => pkt2_0,
          pkt3_0 => pkt3_0,
          pkt4_0 => pkt4_0,
          counter_o => counter_o,
          ethertype_o => ethertype_o,
          ethervalue_o => ethervalue_o,
          counter_index => counter_index,
          grantportint_o => grantportint_o,
          addlpointer_o => addlpointer_o,
          addrpointer_o => addrpointer_o,
          ready2push_o => ready2push_o,
          dropped_o => dropped_o,
          isfull_o => isfull_o,
          clk => clk,
          rst => rst
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '1';
		wait for clk_period/2;
		clk <= '0';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData4 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData5 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData6 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData7 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData8 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData9 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData10 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData11 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData12 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData13 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData14 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData15 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData16 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData17 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData18 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData19 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData20 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData21 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData22 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData23 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData24 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData25 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData26 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData27 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		 iData28 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData29 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData30 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData31 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '1';
       wait for clk_period;

       rst <= '0';
       wait for clk_period*5;


       iData_av <= "00000000000000000000000000000001";
       valid_in <= '0';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period*4;

       iData_av <= "00000000000000000000000000000001";
       iData0 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       valid_in <='1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "0100000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "00001000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;
		 
		  iData_av <= "00000000000000000000000000000000";
       iData0 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '1';
       wait for clk_period;
		 
		 iData_av <= "00000000000000000000000000000001";
		 iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

       valid_in <= '0';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period*15;

       iData_av <= "00000000000000000000000000000001";
       iData0 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       valid_in <='1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "0100000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "00001000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '1';
       wait for clk_period;
		
       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period*8;

       iData_av <= "00000000000000000000000000000100";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;
		 
		 oData_rd <= '0';
		 wait for clk_period*4;

       iData_av <= "00000000000000000000000000000100";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData2 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       valid_in <='1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000010" & "0000000000000011" & "00000010" & "00000000" & "00010000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '1';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData2 <= "00001100000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period*80;

        -- TestCase 2
        -- TestCase 2
        -- TestCase 2
       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period*5;


       iData_av <= "00000000000000000000000000001000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period*4;

       iData_av <= "00000000000000000000000000001000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData3 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00010000" & "0000000000000000";
       valid_in <='1';
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000010000000000" & "0000010000000000" & "00011000" & "00010010" & "10000010" & "00000000" & "00100110" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010111";
       oData_rd <= '0';
       Rd_opcode <= '1';
       rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "00001000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData2 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '1';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       --rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       --rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       --rst <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       wait for clk_period*8;

       iData_av <= "00000000000000000000000000000010";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000010";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData2 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       valid_in <='1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0100000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '1';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       iData2 <= "00001100000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period;

       iData_av <= "00000000000000000000000000000000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid_in <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       wait for clk_period*80;
      wait;
   end process;

END;
