LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY classify_tb IS
END classify_tb;

ARCHITECTURE behavior OF classify_tb IS

    COMPONENT classify_packet
    PORT(
           iData_av : in  STD_LOGIC_VECTOR (3 downto 0);
           iRd_Data : out  STD_LOGIC_VECTOR (3 downto 0);
           iData0 : in  STD_LOGIC_VECTOR (143 downto 0);
           iData1 : in  STD_LOGIC_VECTOR (143 downto 0);
           iData2 : in  STD_LOGIC_VECTOR (143 downto 0);
           iData3 : in  STD_LOGIC_VECTOR (143 downto 0);
           oData_av : out  STD_LOGIC;
           oData_rd : in STD_LOGIC;
           oData : out  STD_LOGIC_VECTOR (143 downto 0);
           MAC : in  STD_LOGIC_VECTOR(47 downto 0);
           valid : in STD_LOGIC;
           Opcode : out  STD_LOGIC_VECTOR(2 downto 0);
           Rd_opcode : in  STD_LOGIC;
           Input_port : out  STD_LOGIC_VECTOR (3 downto 0);
           Port_mask : out  STD_LOGIC_VECTOR (3 downto 0);
           Edge_ports : inout  STD_LOGIC_VECTOR (3 downto 0);
           Core_Ports : inout  STD_LOGIC_VECTOR (3 downto 0);
           gport : out  STD_LOGIC_VECTOR (3 downto 0);  --debug
           ostatus : out STD_LOGIC_VECTOR(1 downto 0); --debug
           oreadstatus : out STD_LOGIC_VECTOR(3 downto 0); --debug
           debug : inout STD_LOGIC_VECTOR(1 downto 0); --debug
           hoppointer_o : out STD_LOGIC_VECTOR(1 downto 0); --debug
           pkt0_0 : out STD_LOGIC_VECTOR(143 downto 0);  --debug
           pkt1_0 : out STD_LOGIC_VECTOR(143 downto 0);  --debug
           pkt2_0 : out STD_LOGIC_VECTOR(143 downto 0);  --debug
           pkt3_0 : out STD_LOGIC_VECTOR(143 downto 0);  --debug
           pkt4_0 : out STD_LOGIC_VECTOR(143 downto 0);  --debug
           counter_o : out STD_LOGIC_VECTOR(3 downto 0); --debug
           ethertype_o : out STD_LOGIC; --debug
           ethervalue_o : out STD_LOGIC; --debug
           counter_index : out integer range 0 to 15; --debug
           grantportint_o : out integer range 1 to 4;   --debug
           addlpointer_o : out integer range 1 to 4;   --debug
           addrpointer_o : out integer range 1 to 4;   --debug
           clk : in  STD_LOGIC;
           rst : in  STD_LOGIC
        );
    END COMPONENT;
    
   --Inputs
   signal iData_av : std_logic_vector(3 downto 0) := (others => '0');
   signal iData0 : std_logic_vector(143 downto 0) := (others => '0');
   signal iData1 : std_logic_vector(143 downto 0) := (others => '0');
   signal iData2 : std_logic_vector(143 downto 0) := (others => '0');
   signal iData3 : std_logic_vector(143 downto 0) := (others => '0');
   signal MAC : std_logic_vector(47 downto 0) := (others => '0');
   signal valid : std_logic := '0';
   signal Rd_opcode : std_logic := '0';
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal oData_rd : STD_LOGIC;

   --Outputs
   signal iRd_Data : std_logic_vector(3 downto 0);
   signal oData_av : std_logic;
   signal oData : std_logic_vector(143 downto 0);
   signal Opcode : std_logic_vector(2 downto 0);
   signal Input_port : std_logic_vector(3 downto 0);
   signal Port_mask : std_logic_vector(3 downto 0);
   signal Edge_ports : std_logic_vector(3 downto 0);
   signal Core_Ports : std_logic_vector(3 downto 0);
   signal gport : STD_LOGIC_VECTOR (3 downto 0);  --debug
   signal ostatus : STD_LOGIC_VECTOR(1 downto 0); --debug
   signal oreadstatus : STD_LOGIC_VECTOR(3 downto 0); --debug
   signal debug : STD_LOGIC_VECTOR(1 downto 0); --debug
   signal hoppointer_o : STD_LOGIC_VECTOR(1 downto 0); --debug
   signal pkt0_0 : STD_LOGIC_VECTOR(143 downto 0);  --debug
   signal pkt1_0 : STD_LOGIC_VECTOR(143 downto 0);  --debug
   signal pkt2_0 : STD_LOGIC_VECTOR(143 downto 0);  --debug
   signal pkt3_0 : STD_LOGIC_VECTOR(143 downto 0);  --debug
   signal pkt4_0 : STD_LOGIC_VECTOR(143 downto 0);  --debug
   signal counter_o : STD_LOGIC_VECTOR(3 downto 0); --debug;
   signal ethertype_o : STD_LOGIC; --debug
   signal ethervalue_o : STD_LOGIC; --debug
   signal counter_index : integer range 0 to 15; --debug
   signal grantportint_o : integer range 1 to 4;   --debug
   signal addlpointer_o : integer range 1 to 4;   --debug
   signal addrpointer_o : integer range 1 to 4;   --debug

   -- Clock period definitions
   constant clk_period : time := 100 ns;

BEGIN

    -- Instantiate the Unit Under Test (UUT)
   uut: classify_packet PORT MAP (
          iData_av => iData_av,
          iRd_Data => iRd_Data,
          iData0 => iData0,
          iData1 => iData1,
          iData2 => iData2,
          iData3 => iData3,
          oData_av => oData_av,
          oData_rd => oData_rd,
          oData => oData,
          MAC => MAC,
          valid => valid,
          Opcode => Opcode,
          Rd_opcode => Rd_opcode,
          Input_port => Input_port,
          Port_mask => Port_mask,
          Edge_ports => Edge_ports,
          Core_Ports => Core_Ports,
          gport => gport,  --debug
          ostatus => ostatus, --debug
          oreadstatus => oreadstatus, --debug
          debug => debug, --debug
          hoppointer_o => hoppointer_o, --debug
          pkt0_0 => pkt0_0, --debug
          pkt1_0 => pkt1_0, --debug
          pkt2_0 => pkt2_0, --debug
          pkt3_0 => pkt3_0, --debug
          pkt4_0 => pkt4_0, --debug
          counter_o => counter_o, --debug
          ethertype_o => ethertype_o,  --debug
          ethervalue_o => ethervalue_o,  --debug
          counter_index => counter_index,  --debug
          grantportint_o => grantportint_o,  --debug
          addlpointer_o => addlpointer_o, --debug
          addrpointer_o => addrpointer_o,  --debug
          clk => clk,
          rst => rst
        );

   -- Clock process definitions
   clk_process :process
   begin
       clk <= '1';
       wait for clk_period/2;
       clk <= '0';
       wait for clk_period/2;
   end process;

   -- Stimulus process
   stim_proc: process
   begin
      -- hold reset state for 100 ns.

      -- insert stimulus here
        -- TestCase 1
       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '1';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*5;


       iData_av <= "0001";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0001";
       iData0 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       valid <='1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "0100000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '1';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "00001000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData2 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*8;

       iData_av <= "0100";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0100";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData2 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       valid <='1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0100000000001010" & "0000000000000011" & "00000010" & "00000000" & "00010000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '1';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData2 <= "00001100000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*80;

        -- TestCase 2
        -- TestCase 2
        -- TestCase 2
       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '1';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*5;


       iData_av <= "1000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "1000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData3 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00010000" & "0000000000000000";
       valid <='1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0100000000000000" & "0000010000000000" & "00011000" & "00010010" & "10000010" & "00000000" & "00100110" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '1';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "00001000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData2 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '0';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*8;

       iData_av <= "0010";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0010";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000001" & "0000000000000000";
       iData2 <= "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "00000000" & "0000000000000000";
       valid <='1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData1 <= "0100000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData2 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       iData3 <= "0000000000000000" & "0000000000000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '1';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "010101010101010101010101010101010101010101010101" & "0000000000000000";
       iData2 <= "00001100000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       iData3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000" & "000000000000000000000000000000000000000000000000" & "0000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '1';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period;

       iData_av <= "0000";
       iData0 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData1 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData2 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       iData3 <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
       valid <= '0';
       MAC <= "010101010101010101010101010101010101010101010101";
       oData_rd <= '1';
       Rd_opcode <= '0';
       rst <= '0';
       wait for clk_period*80;
      wait;
   end process;

END;
